----------------------------------------------------------
--! @file alu_tb
--! @A alu_tb can combine multipal counter to count.
-- Filename: alu_tb.vhd
-- Description: A alu_tb can test the reaction of a register file.
-- Author: YIN Haoping
-- Date: March 27, 2023
----------------------------------------------------------
--! Use standard library
LIBRARY ieee;
use ieee.std_logic_1164.all;
USE ieee.numeric_std.ALL;

--! alu_pkg package description

--! Detailed description of this
--! alu_pkg design element.
PACKAGE alu_pkg IS
--! alu_pkg package description

--! Detailed description of this
--! alu_pkg design element.
	constant ALU_ADD : std_logic_vector(3 downto 0) := "0000";
	constant ALU_SUB : std_logic_vector(3 downto 0) := "0001";
	constant ALU_SLL : std_logic_vector(3 downto 0) := "0010";
	constant ALU_SRL : std_logic_vector(3 downto 0) := "0011";
	constant ALU_SRA : std_logic_vector(3 downto 0) := "0100";
	constant ALU_AND : std_logic_vector(3 downto 0) := "0101";
	constant ALU_OR  : std_logic_vector(3 downto 0) := "0110";
	constant ALU_XOR : std_logic_vector(3 downto 0) := "0111";
	constant ALU_BEQ : std_logic_vector(3 downto 0) := "1000";
	constant ALU_BLT : std_logic_vector(3 downto 0) := "1001";
	constant ALU_BLTU : std_logic_vector(3 downto 0) := "1010";
	constant ALU_JAL : std_logic_vector(3 downto 0) := "1011";
	constant ALU_LUI : std_logic_vector(3 downto 0) := "1100";

	type test_t is
	record
	  op1                         : std_logic_vector(31 downto 0);
	  op2                         : std_logic_vector(31 downto 0);
	  selop                       : std_logic_vector(3 downto 0);
	  exp_res                     : std_logic_vector(31 downto 0);
	  exp_flags                   : std_logic_vector(2 downto 0); -- (0) is EQ flag, (1) is LT flag, (2) is the LTU flag
	end record;
	type test_vectors_t is array (0 to 96) of test_t;

	CONSTANT vectors: test_vectors_t := (
    -- 							op1                 op2                 		selop    			exp_res             exp_flags
	-- ADD
    ("00000000000000000000000000000001", "00000000000000000000000000000001", ALU_ADD, "00000000000000000000000000000010", "000"), 
	(std_logic_vector(to_unsigned(128, 32)), std_logic_vector(to_unsigned(171, 32)), ALU_ADD, std_logic_vector(to_unsigned(299, 32)), "000"),
	(std_logic_vector(to_unsigned(55, 32)), std_logic_vector(to_unsigned(45, 32)), ALU_ADD, std_logic_vector(to_unsigned(100, 32)), "000"),
	(std_logic_vector(to_unsigned(30, 32)), std_logic_vector(to_unsigned(15, 32)), ALU_ADD, std_logic_vector(to_unsigned(45, 32)), "000"),
	(std_logic_vector(to_unsigned(0, 32)), std_logic_vector(to_unsigned(5, 32)), ALU_ADD, std_logic_vector(to_unsigned(5, 32)), "000"),
	("11111111111111111111111111111111", "11111111111111111111111111111111", ALU_ADD, "11111111111111111111111111111110", "000"), -- ADD(-1 + -1)
	("11111111111111111111111111111111", "00000000000000000000000000000001", ALU_ADD, "00000000000000000000000000000000", "000"), -- ADD(-1 + 1)
	("10000000000000000000000000000000", "10000000000000000000000000000000", ALU_ADD, "00000000000000000000000000000000", "000"), -- ADD(-2147483648 + -2147483648)
	("01111111111111111111111111111111", "00000000000000000000000000000001", ALU_ADD, "10000000000000000000000000000000", "000"), -- ADD(2147483647 + 1) -> Overflow
	("10000000000000000000000000000000", "11111111111111111111111111111111", ALU_ADD, "01111111111111111111111111111111", "000"), -- ADD(-2147483648 + -1) -> Overflow
	("10000000000000000000000000000000", "00000000000000000000000000000000", ALU_ADD, "10000000000000000000000000000000", "000"), -- ADD(-2147483648 + 0)
	("01111111111111111111111111111111", "00000000000000000000000000000000", ALU_ADD, "01111111111111111111111111111111", "000"), -- ADD(2147483647 + 0)
	("00000000000000000000000000000000", "00000000000000000000000000000000", ALU_ADD, "00000000000000000000000000000000", "000"), -- ADD(0 + 0)
	
	-- SUB
    ("00000000000000000000000000000011", "00000000000000000000000000000001", ALU_SUB, "00000000000000000000000000000010", "000"), 
	(std_logic_vector(to_signed(15, 32)), std_logic_vector(to_signed(10, 32)), ALU_SUB, std_logic_vector(to_signed(5, 32)), "000"),
	(std_logic_vector(to_signed(10, 32)), std_logic_vector(to_signed(15, 32)), ALU_SUB, std_logic_vector(to_signed(-5, 32)), "000"),
	(std_logic_vector(to_signed(150, 32)), std_logic_vector(to_signed(149, 32)), ALU_SUB, std_logic_vector(to_signed(1, 32)), "000"),
	(std_logic_vector(to_signed(50, 32)), std_logic_vector(to_signed(110, 32)), ALU_SUB, std_logic_vector(to_signed(-60, 32)), "000"),
	("00000000000000000000000000000010", "00000000000000000000000000000001", ALU_SUB, "00000000000000000000000000000001", "000"), -- SUB(2 - 1)
	("00000000000000000000000000000100", "00000000000000000000000000000010", ALU_SUB, "00000000000000000000000000000010", "000"), -- SUB(4 - 2)
	("11111111111111111111111111111111", "11111111111111111111111111111111", ALU_SUB, "00000000000000000000000000000000", "000"), -- SUB(-1 - -1)
	("11111111111111111111111111111111", "00000000000000000000000000000001", ALU_SUB, "11111111111111111111111111111110", "000"), -- SUB(-1 - 1)
	("10000000000000000000000000000000", "10000000000000000000000000000000", ALU_SUB, "00000000000000000000000000000000", "000"), -- SUB(-2147483648 - -2147483648)
	("01111111111111111111111111111111", "11111111111111111111111111111111", ALU_SUB, "10000000000000000000000000000000", "000"), -- SUB(2147483647 - -1) -> Overflow
	("10000000000000000000000000000000", "00000000000000000000000000000001", ALU_SUB, "01111111111111111111111111111111", "000"), -- SUB(-2147483648 - 1) -> Overflow
	("10000000000000000000000000000000", "00000000000000000000000000000000", ALU_SUB, "10000000000000000000000000000000", "000"), -- SUB(-2147483648 - 0)
	("01111111111111111111111111111111", "00000000000000000000000000000000", ALU_SUB, "01111111111111111111111111111111", "000"), -- SUB(2147483647 - 0)
	("00000000000000000000000000000000", "00000000000000000000000000000000", ALU_SUB, "00000000000000000000000000000000", "000"), -- SUB(0 - 0)
	
	-- SLL
    ("00000000000000000000000000000001", "00000000000000000000000000000001", ALU_SLL, "00000000000000000000000000000010", "000"),
	("00000000000000000000000000000001", "00000000000000000000000000000001", ALU_SLL, "00000000000000000000000000000010", "000"), -- SLL(1 << 1)
	("00000000000000000000000000000001", "00000000000000000000000000000010", ALU_SLL, "00000000000000000000000000000100", "000"), -- SLL(1 << 2)
	("10000000000000000000000000000000", "00000000000000000000000000000001", ALU_SLL, "00000000000000000000000000000000", "000"), -- SLL(-2147483648 << 1)
	("01111111111111111111111111111111", "00000000000000000000000000000001", ALU_SLL, "11111111111111111111111111111110", "000"), -- SLL(2147483647 << 1)
	("00000000000000000000000000000000", "00000000000000000000000000000001", ALU_SLL, "00000000000000000000000000000000", "000"), -- SLL(0 << 1)
	("00000000000000000000000000000001", "00000000000000000000000000000000", ALU_SLL, "00000000000000000000000000000001", "000"), -- SLL(1 << 0)
	("00000000000000000000000000000001", "00000000000000000000000000011111", ALU_SLL, "10000000000000000000000000000000", "000"), -- SLL(1 << 31)
	("00000000000000000000000000000010", "00000000000000000000000000011111", ALU_SLL, "00000000000000000000000000000000", "000"), -- SLL(2 << 31)
	
	-- SRL
    ("00000000000000000000000000000010", "00000000000000000000000000000001", ALU_SRL, "00000000000000000000000000000001", "000"), 
	("00000000000000000000000000000010", "00000000000000000000000000000001", ALU_SRL, "00000000000000000000000000000001", "000"), -- SRL(2 >> 1)
	("00000000000000000000000000000100", "00000000000000000000000000000010", ALU_SRL, "00000000000000000000000000000001", "000"), -- SRL(4 >> 2)
	("10000000000000000000000000000000", "00000000000000000000000000000001", ALU_SRL, "01000000000000000000000000000000", "000"), -- SRL(-2147483648 >> 1)
	("01111111111111111111111111111111", "00000000000000000000000000000001", ALU_SRL, "00111111111111111111111111111111", "000"), -- SRL(2147483647 >> 1)
	("00000000000000000000000000000000", "00000000000000000000000000000001", ALU_SRL, "00000000000000000000000000000000", "000"), -- SRL(0 >> 1)
	("00000000000000000000000000000001", "00000000000000000000000000000000", ALU_SRL, "00000000000000000000000000000001", "000"), -- SRL(1 >> 0)
	("10000000000000000000000000000000", "00000000000000000000000000011111", ALU_SRL, "00000000000000000000000000000001", "000"), -- SRL(-2147483648 >> 31)
	("01111111111111111111111111111111", "00000000000000000000000000011111", ALU_SRL, "00000000000000000000000000000000", "000"), -- SRL(2147483647 >> 31)
	
	-- SRA
    ("11111111111111111111111111111110", "00000000000000000000000000000001", ALU_SRA, "11111111111111111111111111111111", "000"), 
	("00000000000000000000000000000010", "00000000000000000000000000000001", ALU_SRA, "00000000000000000000000000000001", "000"), -- SRA(2 >> 1)
	("00000000000000000000000000000100", "00000000000000000000000000000010", ALU_SRA, "00000000000000000000000000000001", "000"), -- SRA(4 >> 2)
	("10000000000000000000000000000000", "00000000000000000000000000000001", ALU_SRA, "11000000000000000000000000000000", "000"), -- SRA(-2147483648 >> 1)
	("01111111111111111111111111111111", "00000000000000000000000000000001", ALU_SRA, "00111111111111111111111111111111", "000"), -- SRA(2147483647 >> 1)
	("00000000000000000000000000000000", "00000000000000000000000000000001", ALU_SRA, "00000000000000000000000000000000", "000"), -- SRA(0 >> 1)
	("00000000000000000000000000000001", "00000000000000000000000000000000", ALU_SRA, "00000000000000000000000000000001", "000"), -- SRA(1 >> 0)
	("10000000000000000000000000000000", "00000000000000000000000000011111", ALU_SRA, "11111111111111111111111111111111", "000"), -- SRA(-2147483648 >> 31)
	("01111111111111111111111111111111", "00000000000000000000000000011111", ALU_SRA, "00000000000000000000000000000000", "000"), -- SRA(2147483647 >> 31)
	
	-- AND
    ("00000000000000000000000000000001", "00000000000000000000000000000000", ALU_AND, "00000000000000000000000000000000", "000"), 
	("00000000000000000000000000001111", "00000000000000000000000000000111", ALU_AND, "00000000000000000000000000000111", "000"), -- AND(15 & 7)
	("00000000000000000000000000010101", "00000000000000000000000000011011", ALU_AND, "00000000000000000000000000010001", "000"), -- AND(21 & 27)
	("10000000000000000000000000000000", "00000000000000000000000000000000", ALU_AND, "00000000000000000000000000000000", "000"), -- AND(-2147483648 & 0)
	("01111111111111111111111111111111", "11111111111111111111111111111111", ALU_AND, "01111111111111111111111111111111", "000"), -- AND(2147483647 & -1)
	("00000000000000000000000000000000", "11111111111111111111111111111111", ALU_AND, "00000000000000000000000000000000", "000"), -- AND(0 & -1)
	("00000000000000000000000000000001", "00000000000000000000000000000000", ALU_AND, "00000000000000000000000000000000", "000"), -- AND(1 & 0)
	
	-- OR
    ("00000000000000000000000000000011", "00000000000000000000000000000101", ALU_OR, "00000000000000000000000000000111", "000"), 
	("00000000000000000000000000001111", "00000000000000000000000000000111", ALU_OR, "00000000000000000000000000001111", "000"), -- OR(15 | 7)
	("00000000000000000000000000010101", "00000000000000000000000000011011", ALU_OR, "00000000000000000000000000011111", "000"), -- OR(21 | 27)
	("10000000000000000000000000000000", "00000000000000000000000000000000", ALU_OR, "10000000000000000000000000000000", "000"), -- OR(-2147483648 | 0)
	("01111111111111111111111111111111", "11111111111111111111111111111111", ALU_OR, "11111111111111111111111111111111", "000"), -- OR(2147483647 | -1)
	("00000000000000000000000000000000", "11111111111111111111111111111111", ALU_OR, "11111111111111111111111111111111", "000"), -- OR(0 | -1)
	("00000000000000000000000000000001", "00000000000000000000000000000000", ALU_OR, "00000000000000000000000000000001", "000"), -- OR(1 | 0)
	
	-- XOR
    ("00000000000000000000000000000001", "00000000000000000000000000000001", ALU_XOR, "00000000000000000000000000000000", "000"), 
	("00000000000000000000000000001111", "00000000000000000000000000000111", ALU_XOR, "00000000000000000000000000001000", "000"), -- XOR(15 ^ 7)
	("00000000000000000000000000010101", "00000000000000000000000000011011", ALU_XOR, "00000000000000000000000000001110", "000"), -- XOR(21 ^ 27)
	("10000000000000000000000000000000", "00000000000000000000000000000000", ALU_XOR, "10000000000000000000000000000000", "000"), -- XOR(-2147483648 ^ 0)
	("01111111111111111111111111111111", "11111111111111111111111111111111", ALU_XOR, "10000000000000000000000000000000", "000"), -- XOR(2147483647 ^ -1)
	("00000000000000000000000000000000", "11111111111111111111111111111111", ALU_XOR, "11111111111111111111111111111111", "000"), -- XOR(0 ^ -1)
	("00000000000000000000000000000001", "00000000000000000000000000000000", ALU_XOR, "00000000000000000000000000000001", "000"), -- XOR(1 ^ 0)
	
	-- BEQ
    ("00000000000000000000000000000011", "00000000000000000000000000000011", ALU_BEQ, "00000000000000000000000000000000", "001"), 
	("00000000000000000000000000001111", "00000000000000000000000000001111", ALU_BEQ, "00000000000000000000000000000000", "001"), -- BEQ(15 == 15)
	("10000000000000000000000000000000", "10000000000000000000000000000000", ALU_BEQ, "00000000000000000000000000000000", "001"), -- BEQ(-2147483648 == -2147483648)
	("00000000000000000000000000001111", "00000000000000000000000000000111", ALU_BEQ, "00000000000000000000000000000000", "000"), -- BEQ(15 != 7)
	("01111111111111111111111111111111", "11111111111111111111111111111111", ALU_BEQ, "00000000000000000000000000000000", "000"), -- BEQ(2147483647 != -1)
	
	-- BLT
    ("00000000000000000000000000000001", "00000000000000000000000000000010", ALU_BLT, "00000000000000000000000000000000", "010"), 
	("11111111111111111111111111111111", "00000000000000000000000000000001", ALU_BLT, "00000000000000000000000000000000", "010"), -- BLT(-1 < 1)
	("00000011111111111111111111111111", "11111111111111111111111111111111", ALU_BLT, "00000000000000000000000000000000", "000"), -- BLT()
	--(std_logic_vector(to_signed(2147483647, 32)), std_logic_vector(to_signed(-2147483648, 32)), ALU_BLT, (others => '0'), "000"),
	("00000000000000000000000000001111", "00000000000000000000000000000111", ALU_BLT, "00000000000000000000000000000000", "000"), -- BLT(15 >= 7)
	("11111111111111111111111111111110", "11111111111111111111111111111111", ALU_BLT, "00000000000000000000000000000000", "010"), -- BLT(-2 < -1)
	
	-- BLTU
	(std_logic_vector(to_unsigned(5, 32)), std_logic_vector(to_unsigned(9, 32)), ALU_BLTU, (others => '0'), "100"),
	("00000000000000000000000000000101", "00000000000000000000000000001001", ALU_BLTU, "00000000000000000000000000000000", "100"), -- BLTU(5 < 9)
	("00000000000000000000000000000001", "00000000000000000000000000001111", ALU_BLTU, "00000000000000000000000000000000", "100"), -- BLTU(1 < 15)
	("00000000000000000000000000001111", "00000000000000000000000000000111", ALU_BLTU, "00000000000000000000000000000000", "000"), -- BLTU(15 >= 7)
	("11111111111111111111111111111110", "11111111111111111111111111111111", ALU_BLTU, "00000000000000000000000000000000", "100"), -- BLTU(4294967294 < 4294967295)
	
	-- JAL
	("00000000000000000000000000000100", "00000000000000000000000000000010", ALU_JAL, "00000000000000000000000000000100", "000"), -- JAL(6) 
	("11111111111111111111111111111110", "00000000000000000000000000000010", ALU_JAL, "11111111111111111111111111111110", "000"), -- JAL(-2)
	("00000000000000000000000000000000", "11111111111111111111111111111110", ALU_JAL, "00000000000000000000000000000000", "000"), -- JAL(0)

	-- LUI
	("00000000000000000000000000000000", "00000000000000000000000000000010", ALU_LUI, "00000000000000000000000000000010", "000"), -- LUI(2)
	("00000000000000000000000000000000", "11111111111111111111111111111111", ALU_LUI, "11111111111111111111111111111111", "000"), -- LUI(-1)
	("00000000000000000000000000000000", "00000000000000000000000000000000", ALU_LUI, "00000000000000000000000000000000", "000")  -- LUI(0)

	
);
	
	
			
	--constant vectors : test_vectors_t := (										-- LTU  LT  EQ flags
	--(std_logic(unsigned(0)), std_logic(unsigned(0)), ALU_ADD, std_logic(unsigned(0)), " 0   0   0" ),
	--(std_logic(unsigned(1)), std_logic(unsigned(1)), "0001", std_logic(unsigned(1)),  " 0   0   0" ),
	--(std_logic(unsigned(2)), std_logic(unsigned(2)), "0010", std_logic(unsigned(2)),  " 0   0   0" )
	--); 
	


component alu is
	--generic(selopbits : positive := 4;flagbits : positive := 3);
	port(
	--INPUTS
	op1 : in std_logic_vector(31 downto 0);
	op2 : in std_logic_vector(31 downto 0);
	selop : in std_logic_vector(3 downto 0);
	--OUTPUTS
	res : out std_logic_vector(31 downto 0);
	flags : out std_logic_vector(2 downto 0)
	);
end component;


END PACKAGE alu_pkg;
