----------------------------------------------------------
--! @file alu_pkg
--! @A alu_pkg can combine multipal counter to count.
-- Filename: alu_pkg.vhd
-- Description: A alu_pkg can test the reaction of a register file.
-- Author: YIN Haoping
-- Date: March 27, 2023
----------------------------------------------------------
--! Use standard library
LIBRARY ieee;
use ieee.std_logic_1164.all;
USE ieee.numeric_std.ALL;

--! alu_pkg package description

--! Detailed description of this
--! alu_pkg design element.
PACKAGE alu_pkg IS
--! alu_pkg package description

--! Detailed description of this
--! alu_pkg design element.
	constant ALU_ADD : std_logic_vector(3 downto 0) := "0000";
	constant ALU_SUB : std_logic_vector(3 downto 0) := "0001";
	constant ALU_SLL : std_logic_vector(3 downto 0) := "0010";
	constant ALU_SRL : std_logic_vector(3 downto 0) := "0011";
	constant ALU_SRA : std_logic_vector(3 downto 0) := "0100";
	constant ALU_AND : std_logic_vector(3 downto 0) := "0101";
	constant ALU_OR  : std_logic_vector(3 downto 0) := "0110";
	constant ALU_XOR : std_logic_vector(3 downto 0) := "0111";
	constant ALU_BEQ : std_logic_vector(3 downto 0) := "1000";
	constant ALU_BLT : std_logic_vector(3 downto 0) := "1001";
	constant ALU_BLTU : std_logic_vector(3 downto 0) := "1010";
	constant ALU_JAL : std_logic_vector(3 downto 0) := "1011";
	constant ALU_LUI : std_logic_vector(3 downto 0) := "1100";
	
	function error_event (alu_code : std_logic_vector(3 downto 0) ) return string;
	
	function change_to_string(data : std_logic_vector) return string;
	
	function to_binary_string(slv : std_logic_vector) return string; 
	
	type test_t is
	record
	  op1                         : std_logic_vector(31 downto 0);
	  op2                         : std_logic_vector(31 downto 0);
	  selop                       : std_logic_vector(3 downto 0);
	  exp_res                     : std_logic_vector(31 downto 0);
	  exp_flags                   : std_logic_vector(2 downto 0); -- (0) is EQ flag, (1) is LT flag, (2) is the LTU flag
	end record;
	type test_vectors_t is array (0 to 200) of test_t;

	CONSTANT vectors: test_vectors_t := (					--each selop shall have enough cases, 16 for exemple.
    -- 							op1                 op2                 		selop    			exp_res             exp_flags
	-- ADD
        -- Test case 1: Basic addition
    ("00000000000000000000000000000100", "00000000000000000000000000000010", ALU_ADD, "00000000000000000000000000000110", "000"),
    -- Test case 2: Adding a larger number to a smaller one
    ("00000000000000000000000000000111", "00000000000000000000000000001000", ALU_ADD, "00000000000000000000000000001111", "000"),
    -- Test case 3: Adding the maximum representable value
    ("00000000000000000000000000000000", "11111111111111111111111111111111", ALU_ADD, "11111111111111111111111111111111", "000"),
    -- Test case 4: Adding the minimum representable value
    ("00000000000000000000000000000000", "00000000000000000000000000000001", ALU_ADD, "00000000000000000000000000000001", "000"),
    -- Test case 5: Adding zero
    ("00000000000000000000000000000101", "00000000000000000000000000000000", ALU_ADD, "00000000000000000000000000000101", "000"),
    -- Test case 6: Adding a number to itself
    ("00000000000000000000000000001100", "00000000000000000000000000001100", ALU_ADD, "00000000000000000000000000011000", "000"),
    -- Test case 7: Adding a negative number
    ("00000000000000000000000000000000", "11111111111111111111111111111011", ALU_ADD, "11111111111111111111111111111011", "000"),
    -- Test case 8: Adding a negative number to a positive number
    ("00000000000000000000000000001001", "11111111111111111111111111111001", ALU_ADD, "00000000000000000000000000000010", "000"),
    -- Test case 9: Adding a positive number to a negative number
    ("11111111111111111111111111110101", "00000000000000000000000000000110", ALU_ADD, "11111111111111111111111111111011", "000"),
    -- Test case 10: Adding to a negative number
    ("11111111111111111111111111110101", "00000000000000000000000000000101", ALU_ADD, "11111111111111111111111111111010", "000"),
    -- Test case 11: Adding the maximum negative number
    ("00000000000000000000000000000000", "10000000000000000000000000000000", ALU_ADD, "10000000000000000000000000000000", "000"),
    -- Test case 12: Adding the maximum positive number to a positive number
    ("00000000000000000000000000000011", "01111111111111111111111111111111", ALU_ADD, "10000000000000000000000000000010", "000"),
    -- Test case 13: Adding the maximum positive number to the maximum negative number
    ("10000000000000000000000000000000", "01111111111111111111111111111111", ALU_ADD, "11111111111111111111111111111111", "000"),
    -- Test case 14: Adding a mid-range positive number to a mid-range negative number
    ("11111111100000000000000000000000", "00000000011111111111111111111111", ALU_ADD, "11111111111111111111111111111111", "000"),	
    -- Test case 15: Adding a mid-range negative number to a mid-range positive number
    ("00000000011111111111111111111111", "11111111100000000000000000000000", ALU_ADD, "11111111111111111111111111111111", "000"),
	-- Test case 16: Maximum positive number added to itself (overflow)
	("01111111111111111111111111111111", "01111111111111111111111111111111", ALU_ADD, "11111111111111111111111111111110", "000"), -- Overflow
	-- Test case 17: Maximum negative number added to itself (overflow)
	("10000000000000000000000000000000", "10000000000000000000000000000000", ALU_ADD, "00000000000000000000000000000000", "100"), -- Overflow
	-- Test case 18: Zero added to maximum positive number (no overflow)
	("00000000000000000000000000000000", "01111111111111111111111111111111", ALU_ADD, "01111111111111111111111111111111", "000"), 
	-- Test case 19: Zero added to maximum negative number (no overflow)
	("00000000000000000000000000000000", "10000000000000000000000000000000", ALU_ADD, "10000000000000000000000000000000", "000"),
	-- Test case 20: Maximum negative number added to maximum positive number (no overflow)
	("10000000000000000000000000000000", "01111111111111111111111111111111", ALU_ADD, "11111111111111111111111111111111", "000"), 
	
	
	-- SUB
    -- Test case 1: Basic subtraction
    ("00000000000000000000000000000100", "00000000000000000000000000000010", ALU_SUB, "00000000000000000000000000000010", "000"),
    -- Test case 2: Subtracting a larger number from a smaller one
    ("00000000000000000000000000000111", "00000000000000000000000000001000", ALU_SUB, "11111111111111111111111111111111", "000"),
    -- Test case 3: Subtracting the maximum representable value
    ("00000000000000000000000000000000", "11111111111111111111111111111111", ALU_SUB, "00000000000000000000000000000001", "000"),
    -- Test case 4: Subtracting the minimum representable value
    ("00000000000000000000000000000000", "00000000000000000000000000000001", ALU_SUB, "11111111111111111111111111111111", "000"),
    -- Test case 5: Subtracting zero
    ("00000000000000000000000000000101", "00000000000000000000000000000000", ALU_SUB, "00000000000000000000000000000101", "000"),
    -- Test case 6: Subtracting a number from itself
    ("00000000000000000000000000001100", "00000000000000000000000000001100", ALU_SUB, "00000000000000000000000000000000", "000"),
    -- Test case 7: Subtracting a negative number
    ("00000000000000000000000000000000", "11111111111111111111111111111011", ALU_SUB, "00000000000000000000000000000101", "000"),
    -- Test case 8: Subtracting a negative number from a positive number
    ("00000000000000000000000000001001", "11111111111111111111111111111001", ALU_SUB, "00000000000000000000000000010000", "000"),
    -- Test case 9: Subtracting a positive number from a negative number
    ("11111111111111111111111111110101", "00000000000000000000000000000110", ALU_SUB, "11111111111111111111111111101111", "000"),	
    -- Test case 10: Subtracting from a negative number
    ("11111111111111111111111111110101", "00000000000000000000000000000101", ALU_SUB, "11111111111111111111111111110000", "000"),	
    -- Test case 11: Subtracting the maximum negative number
    ("00000000000000000000000000000000", "10000000000000000000000000000000", ALU_SUB, "10000000000000000000000000000000", "000"),
    -- Test case 12: Subtracting the maximum positive number from a positive number
    ("00000000000000000000000000001010", "01111111111111111111111111111111", ALU_SUB, "10000000000000000000000000001011", "000"),
    -- Test case 13: Subtracting the maximum positive number from the maximum negative number
    ("10000000000000000000000000000000", "01111111111111111111111111111111", ALU_SUB, "00000000000000000000000000000001", "000"),	--**overflow, out of 32bit
    -- Test case 14: Subtracting a mid-range positive number from a mid-range negative number
    ("11111111100000000000000000000000", "00000000011111111111111111111111", ALU_SUB, "11111111000000000000000000000001", "000"),	--**overflow, out of 32bit
    -- Test case 15: Subtracting a mid-range negative number from a mid-range positive number
    ("00000000011111111111111111111111", "11111111100000000000000000000000", ALU_SUB, "00000000111111111111111111111111", "000"),	
	-- Test case 16: Largest positive number - negative number, should wrap around to largest negative number (2,147,483,647-1)
    ("01111111111111111111111111111111", "00000000000000000000000000000001", ALU_SUB, "01111111111111111111111111111110", "000"),	--**overflow
    -- Test case 17: Largest negative number - positive number, should wrap around to largest positive number
    ("10000000000000000000000000000000", "00000000000000000000000000000001", ALU_SUB, "01111111111111111111111111111111", "000"),
    -- Test case 18: Zero - largest negative number, should return largest positive number+1
    ("00000000000000000000000000000000", "10000000000000000000000000000000", ALU_SUB, "01111111111111111111111111111111", "000"),	--error**overflow, out of the positive limite(01111111111111111111111111111111)
    -- Test case 19: Zero - largest positive number, should return largest negative number+1
    ("00000000000000000000000000000000", "01111111111111111111111111111111", ALU_SUB, "10000000000000000000000000000001", "000"),	
	

	
	
	-- SLL
    -- Test case 1: Shifting a basic number by 1 position
    ("00000000000000000000000000000110", "00000000000000000000000000000001", ALU_SLL, "00000000000000000000000000001100", "000"),
    -- Test case 2: Shifting a basic number by 2 positions
    ("00000000000000000000000000000110", "00000000000000000000000000000010", ALU_SLL, "00000000000000000000000000011000", "000"),
    -- Test case 3: Shifting a basic number by 3 positions
    ("00000000000000000000000000000110", "00000000000000000000000000000011", ALU_SLL, "00000000000000000000000000110000", "000"),
    -- Test case 4: Shifting a large number by 1 position
    ("00000000000000100110011001100110", "00000000000000000000000000000001", ALU_SLL, "00000000000001001100110011001100", "000"),
    -- Test case 5: Shifting a large number by 2 positions
    ("00000000000000100110011001100110", "00000000000000000000000000000010", ALU_SLL, "00000000000010011001100110011000", "000"),
    -- Test case 6: Shifting a large number by 3 positions
    ("00000000000000100110011001100110", "00000000000000000000000000000011", ALU_SLL, "00000000000100110011001100110000", "000"),
    -- Test case 7: Shifting a small number by a large number of positions
    ("00000000000000000000000000000011", "00000000000000000000000000010100", ALU_SLL, "00000000001100000000000000000000", "000"),
    -- Test case 8: Shifting a large number by a large number of positions
    ("00000000000000100110011001100110", "00000000000000000000000000010000", ALU_SLL, "01100110011001100000000000000000", "000"),
    -- Test case 9: Shifting by zero positions
    ("00000000000000100110011001100110", "00000000000000000000000000000000", ALU_SLL, "00000000000000100110011001100110", "000"),
    -- Test case 10: Shifting a zero by 1 position
    ("00000000000000000000000000000000", "00000000000000000000000000000001", ALU_SLL, "00000000000000000000000000000000", "000"),
    -- Test case 11: Shifting a zero by a large number of positions
    ("00000000000000000000000000000000", "00000000000000000000000000010000", ALU_SLL, "00000000000000000000000000000000", "000"),
    -- Test case 12: Shifting a negative number
    ("11111111111111111111111111111001", "00000000000000000000000000000010", ALU_SLL, "11111111111111111111111111100100", "000"),
    -- Test case 13: Shifting a negative number by a large number of positions
    ("11111111111111111111111111111001", "00000000000000000000000000010100", ALU_SLL, "11111111100100000000000000000000", "000"),	--error
    -- Test case 14: Shifting a number with the highest bit set
    ("10000000000000000000000000000000", "00000000000000000000000000000001", ALU_SLL, "00000000000000000000000000000000", "000"),
    -- Test case 15: Shifting a number with the highest bit set by a large number of positions
    ("10000000000000000000000000000000", "00000000000000000000000000010000", ALU_SLL, "00000000000000000000000000000000", "000"),
	-- Test case 16: Shift left the largest negative number by 1, should get zero (as the sign bit is shifted out)
    ("10000000000000000000000000000000", "00000000000000000000000000000001", ALU_SLL, "00000000000000000000000000000000", "000"),
    -- Test case 17: Shift left the smallest positive number by 31, should get the largest negative number (as the sign bit is set)
    ("00000000000000000000000000000001", "00000000000000000000000000011111", ALU_SLL, "10000000000000000000000000000000", "000"),	--error
    -- Test case 18: Shift left zero by any number, should get zero
    ("00000000000000000000000000000000", "00000000000000000000000000011111", ALU_SLL, "00000000000000000000000000000000", "000"),
    -- Test case 19: Shift left any number by zero, should get the same number
    ("01100111000011110000111100001111", "00000000000000000000000000000000", ALU_SLL, "01100111000011110000111100001111", "000"),

	-- SRL
    -- Test case 1: Shifting a basic number by 1 position
    ("00000000000000000000000000001100", "00000000000000000000000000000001", ALU_SRL, "00000000000000000000000000000110", "000"),
    -- Test case 2: Shifting a basic number by 2 positions
    ("00000000000000000000000000001100", "00000000000000000000000000000010", ALU_SRL, "00000000000000000000000000000011", "000"),	
    -- Test case 3: Shifting a basic number by 3 positions
    ("00000000000000000000000000001100", "00000000000000000000000000000011", ALU_SRL, "00000000000000000000000000000001", "000"),	
    -- Test case 4: Shifting a large number by 1 position
    ("00000000000001001100110011001100", "00000000000000000000000000000001", ALU_SRL, "00000000000000100110011001100110", "000"),
    -- Test case 5: Shifting a large number by 2 positions
    ("00000000000010011001100110011000", "00000000000000000000000000000010", ALU_SRL, "00000000000000100110011001100110", "000"),	
    -- Test case 6: Shifting a large number by 3 positions
    ("00000000000100110011001100110000", "00000000000000000000000000000011", ALU_SRL, "00000000000000100110011001100110", "000"),	
    -- Test case 7: Shifting a small number by a large number of positions
    ("00000000001100000000000000000000", "00000000000000000000000000010100", ALU_SRL, "00000000000000000000000000000011", "000"),	
    -- Test case 8: Shifting a large number by a large number of positions
    ("01100110011001100000000000000000", "00000000000000000000000000010000", ALU_SRL, "00000000000000000110011001100110", "000"),	
    -- Test case 9: Shifting by zero positions
    ("00000000000000100110011001100110", "00000000000000000000000000000000", ALU_SRL, "00000000000000100110011001100110", "000"),
    -- Test case 10: Shifting a zero by 1 position
    ("00000000000000000000000000000000", "00000000000000000000000000000001", ALU_SRL, "00000000000000000000000000000000", "000"),
    -- Test case 11: Shifting a zero by a large number of positions
    ("00000000000000000000000000000000", "00000000000000000000000000010000", ALU_SRL, "00000000000000000000000000000000", "000"),
    -- Test case 12: Shifting a negative number
    ("11111111111111111111111111111001", "00000000000000000000000000000010", ALU_SRL, "00111111111111111111111111111110", "000"),
    -- Test case 13: Shifting a negative number by a large number of positions
    ("11111111111111111111111111111001", "00000000000000000000000000010100", ALU_SRL, "00000000000000000000111111111111", "000"),	--error
    -- Test case 14: Shifting a number with the highest bit set
    ("10000000000000000000000000000000", "00000000000000000000000000000001", ALU_SRL, "01000000000000000000000000000000", "000"),
    -- Test case 15: Shifting a number with the highest bit set by a large number of positions
    ("10000000000000000000000000000000", "00000000000000000000000000010000", ALU_SRL, "00000000000000001000000000000000", "000"),	--error
	-- Test case 16: Shift right the smallest positive number by 1, should get zero (as the last bit is shifted out)
    ("00000000000000000000000000000001", "00000000000000000000000000000001", ALU_SRL, "00000000000000000000000000000000", "000"),
    -- Test case 17: Shift right the largest negative number by 31, should get the smallest positive number (as the sign bit is shifted out)
    ("10000000000000000000000000000000", "00000000000000000000000000011111", ALU_SRL, "00000000000000000000000000000001", "000"),
    -- Test case 18: Shift right zero by any number, should get zero
    ("00000000000000000000000000000000", "00000000000000000000000000011111", ALU_SRL, "00000000000000000000000000000000", "000"),
    -- Test case 19: Shift right any number by zero, should get the same number
    ("01100111000011110000111100001111", "00000000000000000000000000000000", ALU_SRL, "01100111000011110000111100001111", "000"),


	-- SRA
    -- Test case 1: Shifting a basic number by 1 position
    ("00000000000000000000000000001100", "00000000000000000000000000000001", ALU_SRA, "00000000000000000000000000000110", "000"),
    -- Test case 2: Shifting a basic number by 2 positions
    ("00000000000000000000000000001100", "00000000000000000000000000000010", ALU_SRA, "00000000000000000000000000000011", "000"),
    -- Test case 3: Shifting a negative number by 1 position
    ("11111111111111111111111111111001", "00000000000000000000000000000001", ALU_SRA, "11111111111111111111111111111100", "000"),
    -- Test case 4: Shifting a negative number by 2 positions
    ("11111111111111111111111111111001", "00000000000000000000000000000010", ALU_SRA, "11111111111111111111111111111110", "000"),
    -- Test case 5: Shifting a number with the highest bit set
    ("10000000000000000000000000000000", "00000000000000000000000000000001", ALU_SRA, "11000000000000000000000000000000", "000"),
    -- Test case 6: Shifting a negative number by a large number of positions
    ("11111111111111111111111111111001", "00000000000000000000000000010100", ALU_SRA, "11111111111111111111111111111111", "000"),
    -- Test case 7: Shifting a number with the highest bit set by a large number of positions
    ("10000000000000000000000000000000", "00000000000000000000000000010000", ALU_SRA, "11111111111111111000000000000000", "000"),	
    -- Test case 8: Shifting a zero by 1 position
    ("00000000000000000000000000000000", "00000000000000000000000000000001", ALU_SRA, "00000000000000000000000000000000", "000"),
    -- Test case 9: Shifting a zero by a large number of positions
    ("00000000000000000000000000000000", "00000000000000000000000000010000", ALU_SRA, "00000000000000000000000000000000", "000"),
    -- Test case 10: Shifting by zero positions
    ("00000000000000100110011001100110", "00000000000000000000000000000000", ALU_SRA, "00000000000000100110011001100110", "000"),
    -- Test case 11: Shifting a number by the number of positions equivalent to its width
    ("00000000000000000000000000001100", "00000000000000000000000000100000", ALU_SRA, "00000000000000000000000000000000", "000"),	--error (why got 1100?)
    -- Test case 12: Shifting a negative number by the number of positions equivalent to its width
    ("11111111111111111111111111111001", "00000000000000000000000000100000", ALU_SRA, "11111111111111111111111111111111", "000"),	--error (why got -7?)
    -- Test case 13: Shifting a number with the highest bit set by the number of positions equivalent to its width
    ("10000000000000000000000000000000", "00000000000000000000000000100000", ALU_SRA, "11111111111111111111111111111111", "000"),	--error	(why negative limit?)
    -- Test case 14: Shifting a number with both positive and negative halves
    ("11111111111111111111111100000000", "00000000000000000000000000001111", ALU_SRA, "11111111111111111111111111111111", "000"),	--error	()
    -- Test case 15: Shifting a number with the highest bit set by a large number of positions
    ("10000000000000000000000000000000", "00000000000000000000000000010011", ALU_SRA, "11111111111111111111000000000000", "000"),	--error**
    -- Test case 16: Shift right the smallest positive number by 1, should get zero (as the last bit is shifted out)
    ("00000000000000000000000000000001", "00000000000000000000000000000001", ALU_SRA, "00000000000000000000000000000000", "000"),
    -- Test case 17: Shift right the largest negative number by 31, should still get the largest negative number (as the sign is preserved)
    ("10000000000000000000000000000000", "00000000000000000000000000011111", ALU_SRA, "11111111111111111111111111111111", "000"),	--error**
    -- Test case 18: Shift right zero by any number, should get zero
    ("00000000000000000000000000000000", "00000000000000000000000000011111", ALU_SRA, "00000000000000000000000000000000", "000"),
    -- Test case 19: Shift right any number by zero, should get the same number
    ("01100111000011110000111100001111", "00000000000000000000000000000000", ALU_SRA, "01100111000011110000111100001111", "000"),
	-- Test case 20: Shift right any number by zero, should get the same number
	("01100111000011110000111100001111", "00000000000000000000000000000000", ALU_SRA, "01100111000011110000111100001111", "000"),
	-- Test case 21: Shifting a number from left to right
    ("10000000000000000000000000000000", "00000000000000000000000000011110", ALU_SRA, "11111111111111111111111111111110", "000"),
	
	-- AND
    -- Test case 1: ANDing two simple numbers
    ("00000000000000000000000000001100", "00000000000000000000000000001010", ALU_AND, "00000000000000000000000000001000", "000"),
    -- Test case 2: ANDing a number with itself
    ("00000000000000000000000000001100", "00000000000000000000000000001100", ALU_AND, "00000000000000000000000000001100", "000"),
    -- Test case 3: ANDing a number with zero
    ("00000000000000000000000000001100", "00000000000000000000000000000000", ALU_AND, "00000000000000000000000000000000", "000"),
    -- Test case 4: ANDing a number with all ones
    ("00000000000000000000000000001100", "11111111111111111111111111111111", ALU_AND, "00000000000000000000000000001100", "000"),
    -- Test case 5: ANDing two different numbers
    ("00000000000000000000000010101010", "00000000000000000000000001010101", ALU_AND, "00000000000000000000000000000000", "000"),
    -- Test case 6: ANDing two identical negative numbers
    ("11111111111111111111111111110110", "11111111111111111111111111110110", ALU_AND, "11111111111111111111111111110110", "000"),
    -- Test case 7: ANDing a negative number and a positive number
    ("11111111111111111111111111110110", "00000000000000000000000000001100", ALU_AND, "00000000000000000000000000000100", "000"),
    -- Test case 8: ANDing a negative number and zero
    ("11111111111111111111111111110110", "00000000000000000000000000000000", ALU_AND, "00000000000000000000000000000000", "000"),
    -- Test case 9: ANDing a negative number and all ones
    ("11111111111111111111111111110110", "11111111111111111111111111111111", ALU_AND, "11111111111111111111111111110110", "000"),
    -- Test case 10: ANDing two different negative numbers
    ("11111111111111111111111110101010", "11111111111111111111111101010101", ALU_AND, "11111111111111111111111100000000", "000"),
    -- Test case 11: ANDing maximum positive and negative numbers
    ("01111111111111111111111111111111", "10000000000000000000000000000000", ALU_AND, "00000000000000000000000000000000", "000"),
    -- Test case 12: ANDing a negative number with itself
    ("11111111111111111111111111111111", "11111111111111111111111111111111", ALU_AND, "11111111111111111111111111111111", "000"),
    -- Test case 13: ANDing a number with inverted version of itself
    ("00000000000000000000000010101010", "11111111111111111111111101010101", ALU_AND, "00000000000000000000000000000000", "000"),
    -- Test case 14: ANDing a number with one less than itself
    ("00000000000000000000000000001100", "00000000000000000000000000001011", ALU_AND, "00000000000000000000000000001000", "000"),
    -- Test case 15: ANDing two random numbers
    ("10101010101010101010101010101010", "01010101010101010101010101010101", ALU_AND, "00000000000000000000000000000000", "000"),
    -- Test case 16: AND with zero, should get zero
    ("01100111000011110000111100001111", "00000000000000000000000000000000", ALU_AND, "00000000000000000000000000000000", "000"),
    -- Test case 17: AND with the largest negative number (all bits are 1), should get the same number
    ("01100111000011110000111100001111", "11111111111111111111111111111111", ALU_AND, "01100111000011110000111100001111", "000"),
    -- Test case 18: AND with the same number, should get the same number
    ("01100111000011110000111100001111", "01100111000011110000111100001111", ALU_AND, "01100111000011110000111100001111", "000"),
    -- Test case 19: AND with its own negation, should get zero
    ("01100111000011110000111100001111", "10011000111100001111000011110000", ALU_AND, "00000000000000000000000000000000", "000"),
	
	
	-- OR
    -- Test case 1: ORing two simple numbers
    ("00000000000000000000000000001100", "00000000000000000000000000001010", ALU_OR, "00000000000000000000000000001110", "000"),
    -- Test case 2: ORing a number with itself
    ("00000000000000000000000000001100", "00000000000000000000000000001100", ALU_OR, "00000000000000000000000000001100", "000"),
    -- Test case 3: ORing a number with zero
    ("00000000000000000000000000001100", "00000000000000000000000000000000", ALU_OR, "00000000000000000000000000001100", "000"),
    -- Test case 4: ORing a number with all ones
    ("00000000000000000000000000001100", "11111111111111111111111111111111", ALU_OR, "11111111111111111111111111111111", "000"),
    -- Test case 5: ORing two different numbers
    ("00000000000000000000000010101010", "00000000000000000000000001010101", ALU_OR, "00000000000000000000000011111111", "000"),
    -- Test case 6: ORing two identical negative numbers
    ("11111111111111111111111111110110", "11111111111111111111111111110110", ALU_OR, "11111111111111111111111111110110", "000"),
    -- Test case 7: ORing a negative number and a positive number
    ("11111111111111111111111111110110", "00000000000000000000000000001100", ALU_OR, "11111111111111111111111111111110", "000"),
    -- Test case 8: ORing a negative number and zero
    ("11111111111111111111111111110110", "00000000000000000000000000000000", ALU_OR, "11111111111111111111111111110110", "000"),
    -- Test case 9: ORing a negative number and all ones
    ("11111111111111111111111111110110", "11111111111111111111111111111111", ALU_OR, "11111111111111111111111111111111", "000"),
    -- Test case 10: ORing two different negative numbers
    ("11111111111111111111111110101010", "11111111111111111111111101010101", ALU_OR, "11111111111111111111111111111111", "000"),
    -- Test case 11: ORing maximum positive and negative numbers
    ("01111111111111111111111111111111", "10000000000000000000000000000000", ALU_OR, "11111111111111111111111111111111", "000"),
    -- Test case 12: ORing a negative number with itself
    ("11111111111111111111111111111111", "11111111111111111111111111111111", ALU_OR, "11111111111111111111111111111111", "000"),
    -- Test case 13: ORing a number with inverted version of itself
    ("00000000000000000000000010101010", "11111111111111111111111101010101", ALU_OR, "11111111111111111111111111111111", "000"),
    -- Test case 14: ORing a number with one less than itself
    ("00000000000000000000000000001100", "00000000000000000000000000001011", ALU_OR, "00000000000000000000000000001111", "000"),
    -- Test case 15: ORing two random numbers
    ("10101010101010101010101010101010", "01010101010101010101010101010101", ALU_OR, "11111111111111111111111111111111", "000"),
    -- Test case 16: OR with zero, should get the same number
    ("01100111000011110000111100001111", "00000000000000000000000000000000", ALU_OR, "01100111000011110000111100001111", "000"),
    -- Test case 17: OR with the largest negative number (all bits are 1), should get the largest negative number
    ("01100111000011110000111100001111", "11111111111111111111111111111111", ALU_OR, "11111111111111111111111111111111", "000"),
    -- Test case 18: OR with the same number, should get the same number
    ("01100111000011110000111100001111", "01100111000011110000111100001111", ALU_OR, "01100111000011110000111100001111", "000"),
    -- Test case 19: OR with its own negation, should get the largest negative number
    ("01100111000011110000111100001111", "10011000111100001111000011110000", ALU_OR, "11111111111111111111111111111111", "000"),
	
	-- XOR
    -- Test case 1: XOR with zero, should get the same number
    ("01100111000011110000111100001111", "00000000000000000000000000000000", ALU_XOR, "01100111000011110000111100001111", "000"),
    -- Test case 2: XOR with the largest negative number (all bits are 1), should get the number's negation
    ("01100111000011110000111100001111", "11111111111111111111111111111111", ALU_XOR, "10011000111100001111000011110000", "000"),
    -- Test case 3: XOR with the same number, should get zero
    ("01100111000011110000111100001111", "01100111000011110000111100001111", ALU_XOR, "00000000000000000000000000000000", "000"),
    -- Test case 4: XOR with its own negation, should get the largest negative number
    ("01100111000011110000111100001111", "10011000111100001111000011110000", ALU_XOR, "11111111111111111111111111111111", "000"),
    -- Test case 5-6: XOR with a number, then XOR with the same number again, should get the original number
    ("01100111000011110000111100001111", "10101010101010101010101010101010", ALU_XOR, "11001101101001011010010110100101", "000"),
    ("11001101101001011010010110100101", "10101010101010101010101010101010", ALU_XOR, "01100111000011110000111100001111", "000"),	
    -- Test case 7: XOR with random numbers
    ("10101010101010101010101010101010", "11111111111111111111111111111111", ALU_XOR, "01010101010101010101010101010101", "000"),
    -- Test case 8: XOR with random numbers
    ("10101010101010101010101010101010", "00000000000000000000000000000000", ALU_XOR, "10101010101010101010101010101010", "000"),
    -- Test case 9: XOR with random numbers
    ("10101010101010101010101010101010", "10101010101010101010101010101010", ALU_XOR, "00000000000000000000000000000000", "000"),
    -- Test case 10: XOR with random numbers
    ("10101010101010101010101010101010", "01010101010101010101010101010101", ALU_XOR, "11111111111111111111111111111111", "000"),
    -- Test case 11: XOR with random numbers
    ("01010101010101010101010101010101", "11111111111111111111111111111111", ALU_XOR, "10101010101010101010101010101010", "000"),
    -- Test case 12: XOR with random numbers
    ("01010101010101010101010101010101", "00000000000000000000000000000000", ALU_XOR, "01010101010101010101010101010101", "000"),
    -- Test case 13: XOR with random numbers
    ("01010101010101010101010101010101", "10101010101010101010101010101010", ALU_XOR, "11111111111111111111111111111111", "000"),
    -- Test case 14: XOR with random numbers
    ("01010101010101010101010101010101", "01010101010101010101010101010101", ALU_XOR, "00000000000000000000000000000000", "000"),

	-- BEQ
    -- Test case 1: Two zeros, should be equal
    ("00000000000000000000000000000000", "00000000000000000000000000000000", ALU_BEQ, "00000000000000000000000000000000", "001"), -- Decimal: (0, 0) Equal, EQ flag set
    -- Test case 2: Zero and non-zero, should not be equal
    ("00000000000000000000000000000000", "00000000000000000000000000000001", ALU_BEQ, "00000000000000000000000000000000", "000"), -- Decimal: (0, 1) Not Equal, EQ flag not set
    -- Test case 3: Same non-zero numbers, should be equal
    ("00000000000000000000000000000001", "00000000000000000000000000000001", ALU_BEQ, "00000000000000000000000000000000", "001"), -- Decimal: (1, 1) Equal, EQ flag set
    -- Test case 4: Different non-zero numbers, should not be equal
    ("00000000000000000000000000000001", "00000000000000000000000000000010", ALU_BEQ, "00000000000000000000000000000000", "000"), -- Decimal: (1, 2) Not Equal, EQ flag not set
    -- Test case 5: Random numbers
    ("11111111111111111111111111111111", "11111111111111111111111111111111", ALU_BEQ, "00000000000000000000000000000000", "001"), -- Decimal: (-1, -1) Equal, EQ flag set
    -- Test case 6: Random numbers
    ("11111111111111111111111111111111", "00000000000000000000000000000000", ALU_BEQ, "00000000000000000000000000000000", "000"), -- Decimal: (-1, 0) Not Equal, EQ flag not set
    -- Test case 7: Random numbers
    ("10101010101010101010101010101010", "10101010101010101010101010101010", ALU_BEQ, "00000000000000000000000000000000", "001"), -- Decimal: (2863311530, 2863311530) Equal, EQ flag set
    -- Test case 8: Random numbers
    ("10101010101010101010101010101010", "01010101010101010101010101010101", ALU_BEQ, "00000000000000000000000000000000", "000"), -- Decimal: (2863311530, 1431655765) Not Equal, EQ flag not set
    -- Test case 9: Random numbers
    ("10000000000000000000000000000000", "10000000000000000000000000000000", ALU_BEQ, "00000000000000000000000000000000", "001"), -- Decimal: (2147483648, 2147483648) Equal, EQ flag set
    -- Test case 10: Random numbers
    ("10000000000000000000000000000000", "01000000000000000000000000000000", ALU_BEQ, "00000000000000000000000000000000", "000"), -- Decimal: (2147483648, 1073741824) Not Equal, EQ flag not set
    -- Test case 11: Random numbers
    ("00000000000000000000000000000000", "11111111111111111111111111111111", ALU_BEQ, "00000000000000000000000000000000", "000"), -- Decimal: (0, -1) Not Equal, EQ flag not set
    -- Test case 12: Random numbers
    ("11111111111111111111111111111111", "01111111111111111111111111111111", ALU_BEQ, "00000000000000000000000000000000", "000"), -- Decimal: (-1, 2147483647) Not Equal, EQ flag not set
    -- Test case 13: Random numbers
    ("01111111111111111111111111111111", "01111111111111111111111111111111", ALU_BEQ, "00000000000000000000000000000000", "001"), -- Decimal: (2147483647, 2147483647) Equal, EQ flag set
    -- Test case 14: Random numbers
    ("01111111111111111111111111111111", "11111111111111111111111111111111", ALU_BEQ, "00000000000000000000000000000000", "000"), -- Decimal: (2147483647, -1) Not Equal, EQ flag not set
    -- Test case 15: Random numbers
    ("11001100110011001100110011001100", "11001100110011001100110011001100", ALU_BEQ, "00000000000000000000000000000000", "001"), -- Decimal: (3435973836, 3435973836) Equal, EQ flag set
    -- Test case 16: Random numbers
    ("11001100110011001100110011001100", "00110011001100110011001100110011", ALU_BEQ, "00000000000000000000000000000000", "000"), -- Decimal: (3435973836, 858993459) Not Equal, EQ flag not set
    -- Test case 17: Random numbers
    ("00110011001100110011001100110011", "00110011001100110011001100110011", ALU_BEQ, "00000000000000000000000000000000", "001"), -- Decimal: (858993459, 858993459) Equal, EQ flag set
    -- Test case 18: Random numbers
    ("00110011001100110011001100110011", "11001100110011001100110011001100", ALU_BEQ, "00000000000000000000000000000000", "000"), -- Decimal: (858993459, 3435973836) Not Equal, EQ flag not set

	-- BLT
    -- Test case 1: Two zeros, should not be less than
    ("00000000000000000000000000000000", "00000000000000000000000000000000", ALU_BLT, "00000000000000000000000000000000", "000"), -- Decimal: (0, 0) Not Less Than, LT flag not set
    -- Test case 2: Zero and non-zero, should be less than
    ("00000000000000000000000000000000", "00000000000000000000000000000001", ALU_BLT, "00000000000000000000000000000000", "010"), -- Decimal: (0, 1) Less Than, LT flag set
    -- Test case 3: Same non-zero numbers, should not be less than
    ("00000000000000000000000000000001", "00000000000000000000000000000001", ALU_BLT, "00000000000000000000000000000000", "000"), -- Decimal: (1, 1) Not Less Than, LT flag not set
    -- Test case 4: op1 less than op2, should be less than
    ("00000000000000000000000000000001", "00000000000000000000000000000010", ALU_BLT, "00000000000000000000000000000000", "010"), -- Decimal: (1, 2) Less Than, LT flag set
    -- Test case 5: op1 equal to op2, should not be less than
    ("11111111111111111111111111111111", "11111111111111111111111111111111", ALU_BLT, "00000000000000000000000000000000", "000"), -- Decimal: (-1, -1) Not Less Than, LT flag not set
    -- Test case 6: op1 greater than op2, should not be less than		--error
    ("11111111111111111111111111111111", "00000000000000000000000000000000", ALU_BLT, "00000000000000000000000000000000", "010"), -- Decimal: (-1, 0) Less Than, LT flag set
    -- Test case 7: op1 less than op2, should be less than				--error
    ("10101010101010101010101010101010", "11111111111111111111111111111111", ALU_BLT, "00000000000000000000000000000000", "010"), -- Decimal: (-1431655766, -1) Less Than, LT flag not set
    -- Test case 8: op1 equal to op2, should not be less than
    ("10101010101010101010101010101010", "10101010101010101010101010101010", ALU_BLT, "00000000000000000000000000000000", "000"), -- Decimal: (-1431655766, -1431655766) Not Less Than, LT flag not set
    -- Test case 9: op1 greater than op2, should not be less than		--error
    ("11111111111111111111111111111111", "10101010101010101010101010101010", ALU_BLT, "00000000000000000000000000000000", "000"), -- Decimal: (-1, -1431655766) Not Less Than, LT flag not set
    -- Test case 10: Large numbers, op1 less than op2, should be less than
    ("11100001111000011110000111100001", "11111111111111111111111111111111", ALU_BLT, "00000000000000000000000000000000", "010"), -- Decimal: (-416074956, -1) Less Than, LT flag set
    -- Test case 11: Large numbers, op1 equal to op2, should not be less than
    ("11100001111000011110000111100001", "11100001111000011110000111100001", ALU_BLT, "00000000000000000000000000000000", "000"), -- Decimal: (-416074956, -416074956) Not Less Than, LT flag not set
    -- Test case 12: Large numbers, op1 greater than op2, should not be less than
    ("11111111111111111111111111111111", "11100001111000011110000111100001", ALU_BLT, "00000000000000000000000000000000", "000"), -- Decimal: (-1, -416074956) Not Less Than, LT flag not set
	
	-- BLTU
    -- Test case 1: Two zeros, should not be less than
    ("00000000000000000000000000000000", "00000000000000000000000000000000", ALU_BLTU, "00000000000000000000000000000000", "000"), -- Decimal: (0, 0) Not Less Than, LTU flag not set
    -- Test case 2: Zero and non-zero, should be less than
    ("00000000000000000000000000000000", "00000000000000000000000000000001", ALU_BLTU, "00000000000000000000000000000000", "100"), -- Decimal: (0, 1) Less Than, LTU flag set
    -- Test case 3: Same non-zero numbers, should not be less than
    ("00000000000000000000000000000001", "00000000000000000000000000000001", ALU_BLTU, "00000000000000000000000000000000", "000"), -- Decimal: (1, 1) Not Less Than, LTU flag not set
    -- Test case 4: op1 less than op2, should be less than
    ("00000000000000000000000000000001", "00000000000000000000000000000010", ALU_BLTU, "00000000000000000000000000000000", "100"), -- Decimal: (1, 2) Less Than, LTU flag set
    -- Test case 5: op1 equal to op2, should not be less than
    ("11111111111111111111111111111111", "11111111111111111111111111111111", ALU_BLTU, "00000000000000000000000000000000", "000"), -- Decimal: (4294967295, 4294967295) Not Less Than, LTU flag not set
    -- *Test case 6: op1 greater than op2, should not be less than		
    ("11111111111111111111111111111111", "00000000000000000000000000000000", ALU_BLTU, "00000000000000000000000000000000", "000"), -- Decimal: (4294967295, 0) Not Less Than, LTU flag not set
    -- Test case 7: op1 less than op2, should be less than				
    ("10101010101010101010101010101010", "11111111111111111111111111111111", ALU_BLTU, "00000000000000000000000000000000", "100"), -- Decimal: (2863311530, 4294967295) Less Than, LTU flag set
    -- Test case 8: op1 equal to op2, should not be less than
    ("10101010101010101010101010101010", "10101010101010101010101010101010", ALU_BLTU, "00000000000000000000000000000000", "000"), -- Decimal: (2863311530, 2863311530) Not Less Than, LTU flag not set
    -- Test case 9: op1 greater than op2, should not be less than
    ("11111111111111111111111111111111", "10101010101010101010101010101010", ALU_BLTU, "00000000000000000000000000000000", "000"), -- Decimal: (4294967295, 2863311530) Not Less Than, LTU flag not set
    -- *Test case 10: op1 less than op2, should be less than				
    ("00001111000011110000111100001111", "11110000111100001111000011110000", ALU_BLTU, "00000000000000000000000000000000", "100"), -- Decimal: (404232216, 4042322160) Less Than, LTU flag set
    -- Test case 11: op1 equal to op2, should not be less than			
    ("00001111000011110000111100001111", "00001111000011110000111100001111", ALU_BLTU, "00000000000000000000000000000000", "000"), -- Decimal: (404232216, 404232216) Not Less Than, LTU flag not set
    -- *Test case 12: op1 greater than op2, should not be less than		
    ("11110000111100001111000011110000", "00001111000011110000111100001111", ALU_BLTU, "00000000000000000000000000000000", "000"), -- Decimal: (4042322160, 404232216) Not Less Than, LTU flag not set
    -- Test case 13: Large numbers, op1 less than op2, should be less than		
    ("11100001111000011110000111100001", "11111111111111111111111111111111", ALU_BLTU, "00000000000000000000000000000000", "100"), -- Decimal: (3879731361, 4294967295) Less Than, LTU flag set
    -- Test case 14: Large numbers, op1 equal to op2, should not be less than
    ("11100001111000011110000111100001", "11100001111000011110000111100001", ALU_BLTU, "00000000000000000000000000000000", "000"), -- Decimal: (3879731361, 3879731361) Not Less Than, LTU flag not set
    -- Test case 15: Large numbers, op1 greater than op2, should not be less than
    ("11111111111111111111111111111111", "11100001111000011110000111100001", ALU_BLTU, "00000000000000000000000000000000", "000"),  -- Decimal: (4294967295, 3879731361) Not Less Than, LTU flag not set

	-- JAL
	("00000000000000000000000000000100", "00000000000000000000000000000010", ALU_JAL, "00000000000000000000000000000100", "000"), -- JAL(6) 
	("11111111111111111111111111111110", "00000000000000000000000000000010", ALU_JAL, "11111111111111111111111111111110", "000"), -- JAL(-2)
	("00000000000000000000000000000000", "11111111111111111111111111111110", ALU_JAL, "00000000000000000000000000000000", "000"), -- JAL(0)

	-- LUI
	("00000000000000000000000000000000", "00000000000000000000000000000010", ALU_LUI, "00000000000000000000000000000010", "000"), -- LUI(2)
	("00000000000000000000000000000000", "11111111111111111111111111111111", ALU_LUI, "11111111111111111111111111111111", "000"), -- LUI(-1)
	("00000000000000000000000000000000", "00000000000000000000000000000000", ALU_LUI, "00000000000000000000000000000000", "000")  -- LUI(0)

);
	
	
			
	--constant vectors : test_vectors_t := (										-- LTU  LT  EQ flags
	--(std_logic(unsigned(0)), std_logic(unsigned(0)), ALU_ADD, std_logic(unsigned(0)), " 0   0   0" ),
	--(std_logic(unsigned(1)), std_logic(unsigned(1)), "0001", std_logic(unsigned(1)),  " 0   0   0" ),
	--(std_logic(unsigned(2)), std_logic(unsigned(2)), "0010", std_logic(unsigned(2)),  " 0   0   0" )
	--); 
	


component alu is
	--generic(selopbits : positive := 4;flagbits : positive := 3);
	port(
	--INPUTS
	op1 : in std_logic_vector(31 downto 0);
	op2 : in std_logic_vector(31 downto 0);
	selop : in std_logic_vector(3 downto 0);
	--OUTPUTS
	res : out std_logic_vector(31 downto 0);
	flags : out std_logic_vector(2 downto 0)
	);
end component;


END PACKAGE alu_pkg;


PACKAGE BODY alu_pkg IS

	function change_to_string(data : std_logic_vector) return string is
	begin
		return integer'image(to_integer(unsigned(data)));
	end function change_to_string;

	function error_event (alu_code : std_logic_vector(3 downto 0) ) return string is
	begin
		case alu_code is
			when "0000" =>
				return string'("ALU_ADD");
			when "0001" =>
				return string'("ALU_SUB");
			when "0010" =>
				return string'("ALU_SLL");
			when "0011" =>
				return string'("ALU_SRL");
			when "0100" =>
				return string'("ALU_SRA");
			when "0101" =>
				return string'("ALU_AND");
			when "0110" =>
				return string'("ALU_OR");
			when "0111" =>
				return string'("ALU_XOR");
			when "1000" =>
				return string'("ALU_BEQ");
			when "1001" =>
				return string'("ALU_BLT");
			when "1010" =>
				return string'("ALU_BLTU");
			when "1011" =>
				return string'("ALU_JAL");
			when "1100" =>
				return string'("ALU_LUI");
			when others =>
				return string'("Wrong ALU code");
		end case;
	end function error_event;
	
	
	function to_binary_string(slv : std_logic_vector) return string is
		variable result : string (1 to 32);
	begin
		for i in slv'range loop
			result(i + 1) := std_logic'image(slv(i))(2);
		end loop;
		return result;
	end function to_binary_string;
	
	
END PACKAGE BODY alu_pkg;
